/*
 * MIG7Mock
 * Mock implementation of MIG7 memory controller for simulation
 */
module MIG7Mock #(
    parameter ADDR_WIDTH = 29,        // Address width is in bytes -> 2^29 = 512MB
    parameter DATA_WIDTH = 256,       // Data width is 256 bits = 32 bytes -> 8 words
    parameter MASK_WIDTH = 32,
    parameter RAM_DEPTH  = 33554432,  // Configurable RAM depth in bytes for simulation (32MB for now)
    parameter LIST       = "memory/mig7mock.list" // Initialization file for RAM
) (
    // System interface
    input  wire                     sys_clk_i,
    input  wire                     sys_rst,
    output wire                     ui_clk,
    output wire                     ui_clk_sync_rst,
    output wire                     init_calib_complete,

    // Application interface
    input  wire [ADDR_WIDTH-1:0]    app_addr,
    input  wire [2:0]               app_cmd,
    input  wire                     app_en,
    output wire                     app_rdy,

    // Write data interface
    input  wire [DATA_WIDTH-1:0]    app_wdf_data,
    input  wire                     app_wdf_end,
    input  wire [MASK_WIDTH-1:0]    app_wdf_mask,
    input  wire                     app_wdf_wren,
    output wire                     app_wdf_rdy,

    // Read data interface
    output wire [DATA_WIDTH-1:0]    app_rd_data,
    output wire                     app_rd_data_end,
    output wire                     app_rd_data_valid,

    // Unused signals (tied off)
    input  wire                     app_sr_req,
    input  wire                     app_ref_req,
    input  wire                     app_zq_req,
    output wire                     app_sr_active,
    output wire                     app_ref_ack,
    output wire                     app_zq_ack
);

// Clock and reset generation
assign ui_clk = sys_clk_i;
assign ui_clk_sync_rst = sys_rst;

// Unused signal tie-offs
assign app_sr_active = 1'b0;
assign app_ref_ack = 1'b0;
assign app_zq_ack = 1'b0;

// State machine parameters
localparam INIT_CYCLES = 50;
localparam READ_CYCLES = 10;
localparam WRITE_CYCLES = 10;

// State definitions
localparam INIT = 3'b000;
localparam IDLE = 3'b001;
localparam WRITE_CMD = 3'b010;
localparam WRITE_DATA = 3'b011;
localparam READ_CMD = 3'b100;
localparam READ_DATA = 3'b101;

// Internal registers
reg [2:0] state = 3'b000;
reg [7:0] cycle_counter = 8'd0;
reg init_complete = 1'b0;
reg app_rdy_reg = 1'b0;
reg app_wdf_rdy_reg = 1'b0;
reg [DATA_WIDTH-1:0] app_rd_data_reg = {DATA_WIDTH{1'b0}};
reg app_rd_data_valid_reg = 1'b0;
reg app_rd_data_end_reg = 1'b0;

// Command and address storage
reg [ADDR_WIDTH-1:0] stored_addr = {ADDR_WIDTH{1'b0}};
reg [2:0] stored_cmd = 3'b000;

// RAM storage - depth is in 256-bit words, so divide byte depth by 32
localparam RAM_WORD_DEPTH = RAM_DEPTH / 32; // Convert byte depth to word depth
reg [DATA_WIDTH-1:0] ram_memory [0:RAM_WORD_DEPTH-1];

// Calculate bit width needed for word address
localparam WORD_ADDR_BITS = $clog2(RAM_WORD_DEPTH);
wire [WORD_ADDR_BITS-1:0] ram_word_addr;

// Convert byte address to word address (divide by 32 since 256 bits = 32 bytes)
// We use stored_addr[ADDR_WIDTH-1:5] because dividing by 32 = right shift by 5 bits
assign ram_word_addr = stored_addr[ADDR_WIDTH-1:5];

// Output assignments
assign init_calib_complete = init_complete;
assign app_rdy = app_rdy_reg;
assign app_wdf_rdy = app_wdf_rdy_reg;
assign app_rd_data = app_rd_data_valid_reg ? app_rd_data_reg : {DATA_WIDTH{1'b0}};
assign app_rd_data_valid = app_rd_data_valid_reg;
assign app_rd_data_end = app_rd_data_end_reg;

// Initialize RAM from file
initial begin
    $readmemb(LIST, ram_memory);
end

// Main state machine
always @(posedge ui_clk) begin
    if (ui_clk_sync_rst) begin
        state <= INIT;
        cycle_counter <= 8'd0;
        init_complete <= 1'b0;
        app_rdy_reg <= 1'b0;
        app_wdf_rdy_reg <= 1'b0;
        app_rd_data_reg <= {DATA_WIDTH{1'b0}};
        app_rd_data_valid_reg <= 1'b0;
        app_rd_data_end_reg <= 1'b0;
        stored_addr <= {ADDR_WIDTH{1'b0}};
        stored_cmd <= 3'b000;
    end
    else begin
        case (state)
            INIT: begin
                // Initialization phase
                app_rdy_reg <= 1'b0;
                app_wdf_rdy_reg <= 1'b0;
                app_rd_data_valid_reg <= 1'b0;
                app_rd_data_end_reg <= 1'b0;
                
                if (cycle_counter < INIT_CYCLES - 1) begin
                    cycle_counter <= cycle_counter + 1;
                end
                else begin
                    init_complete <= 1'b1;
                    state <= IDLE;
                    cycle_counter <= 8'd0;
                end
            end
            
            IDLE: begin
                // Ready to accept commands
                app_rdy_reg <= 1'b1;
                app_wdf_rdy_reg <= 1'b1;
                app_rd_data_valid_reg <= 1'b0;
                app_rd_data_end_reg <= 1'b0;
                
                if (app_en && app_rdy_reg) begin
                    stored_addr <= app_addr;
                    stored_cmd <= app_cmd;
                    app_rdy_reg <= 1'b0;
                    cycle_counter <= 8'd0;
                    
                    if (app_cmd == 3'b000) begin // Write command
                        // Check if write data is provided in the same cycle
                        if (app_wdf_wren && app_wdf_rdy_reg && app_wdf_end) begin
                            // Single-cycle write: data is available immediately
                            // Convert byte address to word address for bounds checking
                            if (app_addr < RAM_DEPTH && (app_addr[4:0] == 5'b00000)) begin // Check alignment
                                ram_memory[app_addr[ADDR_WIDTH-1:5]] <= app_wdf_data;
                                $display("%d: MIG7Mock WRITE: byte_addr=0x%h, word_addr=0x%h, data=0x%h", 
                                    $time, app_addr, app_addr[ADDR_WIDTH-1:5], app_wdf_data);
                            end else if (app_addr >= RAM_DEPTH) begin
                                $display("%d: MIG7Mock WRITE OUT-OF-BOUNDS: byte_addr=0x%h (>= 0x%h)", 
                                    $time, app_addr, RAM_DEPTH);
                            end else begin
                                $display("%d: MIG7Mock WRITE UNALIGNED: byte_addr=0x%h (not 32-byte aligned)", 
                                    $time, app_addr);
                            end
                            // Go directly to write processing delay
                            app_wdf_rdy_reg <= 1'b0;
                            state <= WRITE_DATA;
                        end else begin
                            // Multi-cycle write: wait for data in next state
                            state <= WRITE_CMD;
                            app_wdf_rdy_reg <= 1'b1;
                        end
                    end
                    else if (app_cmd == 3'b001) begin // Read command
                        state <= READ_CMD;
                        app_wdf_rdy_reg <= 1'b0;
                    end
                end
            end
            
            WRITE_CMD: begin
                // Wait for write data
                app_rdy_reg <= 1'b0;
                
                if (app_wdf_wren && app_wdf_rdy_reg && app_wdf_end) begin
                    // Write data to RAM (skip mask handling as it will not be used by the design)
                    // Check bounds using byte address and alignment
                    if (stored_addr < RAM_DEPTH && (stored_addr[4:0] == 5'b00000)) begin // Check alignment
                        ram_memory[ram_word_addr] <= app_wdf_data;
                        $display("%d: MIG7Mock WRITE: byte_addr=0x%h, word_addr=0x%h, data=0x%h", 
                            $time, stored_addr, ram_word_addr, app_wdf_data);
                    end else if (stored_addr >= RAM_DEPTH) begin
                        $display("%d: MIG7Mock WRITE OUT-OF-BOUNDS: byte_addr=0x%h (>= 0x%h)", 
                            $time, stored_addr, RAM_DEPTH);
                    end else begin
                        $display("%d: MIG7Mock WRITE UNALIGNED: byte_addr=0x%h (not 32-byte aligned)", 
                            $time, stored_addr);
                    end
                    
                    app_wdf_rdy_reg <= 1'b0;
                    state <= WRITE_DATA;
                    cycle_counter <= 8'd0;
                end
            end
            
            WRITE_DATA: begin
                // Write processing delay
                app_rdy_reg <= 1'b0;
                app_wdf_rdy_reg <= 1'b0;
                
                if (cycle_counter < WRITE_CYCLES - 1) begin
                    cycle_counter <= cycle_counter + 1;
                end
                else begin
                    state <= IDLE;
                    cycle_counter <= 8'd0;
                end
            end
            
            READ_CMD: begin
                // Read processing delay
                app_rdy_reg <= 1'b0;
                app_wdf_rdy_reg <= 1'b0;
                
                if (cycle_counter < READ_CYCLES - 1) begin
                    cycle_counter <= cycle_counter + 1;
                end
                else begin
                    // Load data from RAM
                    // Check bounds using byte address and alignment
                    if (stored_addr < RAM_DEPTH && (stored_addr[4:0] == 5'b00000)) begin // Check alignment
                        app_rd_data_reg <= ram_memory[ram_word_addr];
                        $display("%d: MIG7Mock READ: byte_addr=0x%h, word_addr=0x%h, data=0x%h", 
                            $time, stored_addr, ram_word_addr, ram_memory[ram_word_addr]);
                    end
                    else if (stored_addr >= RAM_DEPTH) begin
                        app_rd_data_reg <= {DATA_WIDTH{1'b0}}; // Return zeros for out-of-bounds
                        $display("%d: MIG7Mock READ OUT-OF-BOUNDS: byte_addr=0x%h (>= 0x%h), returning 0x0", 
                            $time, stored_addr, RAM_DEPTH);
                    end else begin
                        app_rd_data_reg <= {DATA_WIDTH{1'b0}}; // Return zeros for unaligned
                        $display("%d: MIG7Mock READ UNALIGNED: byte_addr=0x%h (not 32-byte aligned), returning 0x0", 
                            $time, stored_addr);
                    end
                    
                    state <= READ_DATA;
                    cycle_counter <= 8'd0;
                end
            end
            
            READ_DATA: begin
                // Output read data
                app_rdy_reg <= 1'b0;
                app_wdf_rdy_reg <= 1'b0;
                app_rd_data_valid_reg <= 1'b1;
                app_rd_data_end_reg <= 1'b1;
                
                // Return to idle after one cycle
                state <= IDLE;
            end
            
            default: begin
                state <= INIT;
            end
        endcase
    end
end

endmodule
